//////////////////////////////////////////////////////////////////////
//          ██╗       ██████╗   ██╗  ██╗    ██████╗            		//
//          ██║       ██╔══█║   ██║  ██║    ██╔══█║            		//
//          ██║       ██████║   ███████║    ██████║            		//
//          ██║       ██╔═══╝   ██╔══██║    ██╔═══╝            		//
//          ███████╗  ██║  	    ██║  ██║    ██║  	           		//
//          ╚══════╝  ╚═╝  	    ╚═╝  ╚═╝    ╚═╝  	           		//
//                                                             		//
// 	2025 Advanced VLSI System Design, Advisor: Lih-Yih, Chiou		//
//                                                             		//
//////////////////////////////////////////////////////////////////////
//                                                             		//
// 	Author: 		                           				  	    //
//	Filename:		top.sv		                                    //
//	Description:	top module for AVSD HW1                     	//
// 	Date:			2025/XX/XX								   		//
// 	Version:		1.0	    								   		//
//////////////////////////////////////////////////////////////////////
`include "SRAM_wrapper.sv"

module top(
input clk,
input rst
);


// --------------------------//
//   Instance Your CPU Here  //
// --------------------------//





SRAM_wrapper IM1(
.CLK(),
.RST(),
.CEB(),
.WEB(),
.BWEB(),
.A(),
.DI(),
.DO()
);

SRAM_wrapper DM1(
.CLK(),
.RST(),
.CEB(),
.WEB(),
.BWEB(),
.A(),
.DI(),
.DO()
);

endmodule